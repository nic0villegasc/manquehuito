`timescale 1ns/1ps

// Copyright 2025 Universidad de los Andes, Chile
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Authors:
// - Nicolás Villegas <navillegas@miuandes.cl>

// -----------------------------------------------------------------------------
// Module: control_unit
// Description: Decodes 7-bit opcode into a 12-bit control signal based on opcode
//              and optionally condition flags (ZNCV).
// -----------------------------------------------------------------------------
module control_unit (
  input  logic [6:0]  opcode_i,  // 7-bit opcode
  input  logic [3:0]  zncv_i,    // Flags: Zero, Negative, Carry, Overflow
  output logic [11:0] out_o      // Decoded control signals
);

  always_comb begin
    out_o = 12'b0;
    unique case (opcode_i)
      'b0000000: out = 12'b000101000000;
      'b0000001: out = 12'b000010011000;
      'b0000010: out = 12'b000101010000;
      'b0000011: out = 12'b000011010000;
      'b0000100: out = 12'b000100000000;
      'b0000101: out = 12'b000010000000;
      'b0000110: out = 12'b000100010000;
      'b0000111: out = 12'b000011110000;
      'b0001000: out = 12'b000100000001;
      'b0001001: out = 12'b000010000001;
      'b0001010: out = 12'b000100010001;
      'b0001011: out = 12'b000011110001;
      'b0001100: out = 12'b000100000010;
      'b0001101: out = 12'b000010000010;
      'b0001110: out = 12'b000100010010;
      'b0001111: out = 12'b000011110010;
      'b0010000: out = 12'b000100000011;
      'b0010001: out = 12'b000010000011;
      'b0010010: out = 12'b000100010011;
      'b0010011: out = 12'b000011110011;
      'b0010100: out = 12'b000100000100;
      'b0010101: out = 12'b000101100100;
      'b0010110: out = 12'b000010000100;
      'b0010111: out = 12'b000011100100;
      'b0011000: out = 12'b000100000101;
      'b0011001: out = 12'b000010000101;
      'b0011010: out = 12'b000100010101;
      'b0011011: out = 12'b000011110101;
      'b0011100: out = 12'b000100000110;
      'b0011101: out = 12'b000101100110;
      'b0011110: out = 12'b000010000110;
      'b0011111: out = 12'b000011100110;
      'b0100000: out = 12'b000100000111;
      'b0100001: out = 12'b000101100111;
      'b0100010: out = 12'b000010000111;
      'b0100011: out = 12'b000011100111;
      'b0100100: out = 12'b000010100000;
      'b0100101: out = 12'b000101001000;
      'b0100110: out = 12'b000011001000;
      'b0100111: out = 12'b010000011000;
      'b0101000: out = 12'b010001000000;
      'b0101001: out = 12'b001101001000;
      'b0101010: out = 12'b001011001000;
      'b0101011: out = 12'b011000011000;
      'b0101100: out = 12'b000100001000;
      'b0101101: out = 12'b000011101000;
      'b0101110: out = 12'b001100001000;
      'b0101111: out = 12'b010000000000;
      'b0110000: out = 12'b000100001001;
      'b0110001: out = 12'b000011101001;
      'b0110010: out = 12'b001100001001;
      'b0110011: out = 12'b010000000001;
      'b0110100: out = 12'b000100001010;
      'b0110101: out = 12'b000011101010;
      'b0110110: out = 12'b001100001010;
      'b0110111: out = 12'b010000000010;
      'b0111000: out = 12'b000100001011;
      'b0111001: out = 12'b000011101011;
      'b0111010: out = 12'b001100001011;
      'b0111011: out = 12'b010000000011;
      'b0111100: out = 12'b010000000100;
      'b0111101: out = 12'b010001100100;
      'b0111110: out = 12'b011000000100;
      'b0111111: out = 12'b000100001101;
      'b1000000: out = 12'b000011101101;
      'b1000001: out = 12'b001100001101;
      'b1000010: out = 12'b010000000101;
      'b1000011: out = 12'b010000000110;
      'b1000100: out = 12'b010001100110;
      'b1000101: out = 12'b011000000110;
      'b1000110: out = 12'b010000000111;
      'b1000111: out = 12'b010001100111;
      'b1001000: out = 12'b011000000111;
      'b1001001: out = 12'b010000101000;
      'b1001010: out = 12'b011000101000;
      'b1001011: out = 12'b010001011000;
      'b1001100: out = 12'b011001011000;
      'b1001101: out = 12'b000000000001;
      'b1001110: out = 12'b000000010001;
      'b1001111: out = 12'b000001110001;
      'b1010000: out = 12'b000000001001;
      'b1010001: out = 12'b000001101001;
      'b1010010: out = 12'b001000001001;
      'b1010011: out = 12'b100000000000;

      7'b1010100: if (zncv_i[3])                   out_o = 12'b100000000000; // Z == 1
      7'b1010101: if (!zncv_i[3])                  out_o = 12'b100000000000; // Z == 0
      7'b1010110: if (!zncv_i[3] && !zncv_i[2])    out_o = 12'b100000000000; // Z == 0 && N == 0
      7'b1010111: if (zncv_i[2])                   out_o = 12'b100000000000; // N == 1
      7'b1011000: if (!zncv_i[2])                  out_o = 12'b100000000000; // N == 0
      7'b1011001: if (zncv_i[3] || zncv_i[2])      out_o = 12'b100000000000; // Z == 1 || N == 1
      7'b1011010: if (zncv_i[1])                   out_o = 12'b100000000000; // C == 1
      7'b1011011: if (zncv_i[0])                   out_o = 12'b100000000000; // V == 1
    endcase
  end

endmodule : control_unit